library ieee;

entity F_Split is
  port( SR_E:   in Bit_vector(23 downto 0);
        clk:    in Bit;
        SR_Fs:  out Bit_vector(23 downto 0);
end F_Split;

architecture frequenzysplit of F_Split is
begin
    --zeuch das frequenz teilt..
    
    
    
end
  


